

module AXI4_SHIFT(
    // AXI4 BUS
    input wire ACLK,
    input wire ARESETn,
    input wire TKEEP,
    input wire TSTRB,
    input wire TDATA
);
    
endmodule